/* Заметки:
1. Для штатной работы однотактного ядра (SINGLECYCLE_CORE) необходима асинхронная память инструкций
и данных, которая может быть получена при варианте синтезируемой на ячейках памяти(SYNTH_MEM). В
таком режиме ядро практически полностью является комбинационным и может работать на общей частоте
тактирования (clk), одна инструкция выполняется за один такт. Если же использовать внутреннюю
память плис (BSRAM_MEM), которая является синхронной, то ядро становистя псевдо однотактным
поскольку данные записываются и считываются из памяти по переднему фронту тактового сигнала и для
одной инструкции необходимо уже 3 такта. Первый такт приходит на тактирования всех узлов ядра,
кроме памяти инструкций, которая тактируется от второго такта, и памяти данных, которая тактируется
от третьего такта. Думаю что реализвация однотактного ядра с синхронной памятью возможна при
2 тактах, необходима !дополнительная проработка!
2. При использовании памяти BSRAM в конвеерном ядре межстадийным регистром является сама память
поскольку она явлется синхронной и выдаёт данные на выход по такту. При использовании синтезированной
памяти в конвеерном ядре нужен дополнительный межстадийный регистр поскольку память асинхронная и
необходимо разделить стадии регистрами. Для однотактного ядра межстадийный регистр не нужен, связь
явлется проводником.
3. Связано с пунктом 2. При разработке приостановки конвейера, всвязи с конфликтом при выполнении
инструкции lw, необходимо задержать межстадийный регистр (fetch-decode) на один такт. Поскольку в
конвейерном ядре с памятью BSRAM межстадийным регистром является сама память приходится отключать
тактирование памяти на 1 такт подачей сигнала imem_re на контакт ce (clock enable) BSRAM. В текущей
конфигурации кода появилось очень длинная связь именно логическая, сложная для понимания, но не
нарушающая и не ухудшающая параметры ядра. Возможно пересмотреть.
4. Не очень нравится как реализованы интерфейсы мамяти в ядре. Может лучше достать их из модулей
стадий конвейера и поместить в главный модуль core. Подумать.
5. Можно сократить одну операцию в модуле АЛУ, если объединить вместе операции арифметического
и логического сдвига с предварительной подготовкой знакового бита, согласно следующему выражению:
3'b111: ALUResult = $signed({($sra | $srai) ? srcA[31] : 1'b0, srcA}) >>> srcB[4:0];
В таком случае также можно будет уменьшить разрядность ALUControl до 3ёх, но потребуется дополнительные
флаги о том что выполняется команда sra или srai.
6. Упёрся в частоту при синтезировании однотактного ядра на этапе добавления блока загрузки/выгрузки (LSU).
Частота процессора 27MHz. А в проблемной конфигурации (однотактное ядро с синтезированной памятью)
частота ещё в 3 раза ниже. Можно немного немного уменьшить временные задержки, если сделать несколько
параллельных цепей расширения знака. Возможно это повлияет на работу конвейерного ядра при увеличении
частоты, необходимо обратить на это внимание в дальнейшем. 
*/

//============================================================================================== 
// Определения настроек ядра
//============================================================================================== 
//#1 CORE_TYPE #
`define SINGLECYCLE_CORE 1
`define PIPELINE_CORE    0
//#2 MEMORY_TYPE #
`define BSRAM_MEM        1
`define SYNTH_MEM        0
//DSECRIPTION:
//1) Максимальная суммарная память BSRAM_IMEM_SIZE + BSRAM_DMEM_SIZE = 48кБ.
//============================================================================================== 
    
module top #(parameter bit CORE_TYPE       = `SINGLECYCLE_CORE,
                //Настройки памяти инструкций
             parameter bit IMEM_TYPE       =        `BSRAM_MEM,
             parameter int BSRAM_IMEM_SIZE =                 8, //кБайт (поддерживаемые значения 8/16/32)
             parameter int SYNTH_IMEM_SIZE =               100, //слов по 4 Байт
             parameter     IMEM_INIT_FILE  =  "mem_init/i.mem",
                //Настройки памяти данных
             parameter bit DMEM_TYPE       =        `BSRAM_MEM,
             parameter int BSRAM_DMEM_SIZE =                 8, //кБайт (поддерживаемые значения 8/16/32)
             parameter int SYNTH_DMEM_SIZE =                10, //слов по 4 Байт
             parameter     DMEM_INIT_FILE  =  "mem_init/d.mem")   
            (input  logic       clk,     //Вход тактирования
             input  logic       rst_n,   //Вход сброса (кнопка S2)
             output logic [5:0] led      //Выход на 6 светодиодов
);
    //#0 Настройка тактирования
    //DESCRIPTION: Для однотактного ядра при использовании BSAM делаем псевдооднотактный процессор
    //с тремя тактами на одну инструкцию. Тактируем imem и dmem 2ым и 3ьим тактом.
    logic clk_div2;
    always_ff @(posedge clk) clk_div2 <= ~clk_div2;

    logic clk_core, clk_imem, clk_dmem;
    generate if ((IMEM_TYPE | DMEM_TYPE) & CORE_TYPE) begin   //#1 - Для однотактного ядра с BSRAM
        divideby3 divideby3(.clk(clk_div2), .clk_div3(clk_core), .clk_imem(clk_imem), .clk_dmem(clk_dmem));
    end else begin                                            //#0 - Прочие конфигурации
        assign clk_core = clk_div2;
        assign clk_imem = clk_div2;
        assign clk_dmem = clk_div2;
    end
    endgenerate
    
    //#1 Устранение дребезжания с кнопки S2 (rst_n)
    logic [15:0] btn_sync = 0;
    logic rst_sync_n = 0;
    logic rst_sync;
    
    always_ff @(posedge clk_core)
        if (rst_n)
            btn_sync <= {btn_sync[14:0], 1'b1};
        else
            btn_sync <= {1'b0, btn_sync[15:1]};
    
    always_ff @(posedge clk_core) 
        if (btn_sync == 16'b1111_1111_1111_1111) rst_sync_n <= 1'b1;
        else    if (btn_sync == 16'b0000_0000_0000_0000) rst_sync_n <= 1'b0;
                else rst_sync_n <= rst_sync_n;

    assign rst_sync = ~rst_sync_n;

    //#2 Подключаем ядро процессора
        //Интерфейс памяти команд
    logic [31:0] imem_data;
    logic        imem_re, imem_rst;
    logic [31:0] imem_addr;
        //Интерфейс памяти данных
    logic [31:0] dmem_ReadData;
    logic [ 3:0] dmem_Write;
    logic [31:0] dmem_Addr, dmem_WriteData;
        //Ядро
    core #(CORE_TYPE, IMEM_TYPE, DMEM_TYPE)
           riscv  
          (.clk(clk_core), .rst(rst_sync), .out(led),                                            //Системные
           .imem_data(imem_data), .imem_re(imem_re), .imem_rst(imem_rst), .imem_addr(imem_addr), //Интерфейс памяти команд
           .dmem_ReadData(dmem_ReadData), .dmem_Write(dmem_Write),                               //Интерфейс памяти данных
           .dmem_Addr(dmem_Addr), .dmem_WriteData(dmem_WriteData));
   
    //#3 Подключаем память
    mem #(IMEM_TYPE, SYNTH_IMEM_SIZE, BSRAM_IMEM_SIZE, IMEM_INIT_FILE) imem
          (.clk(clk_imem), .reset(rst_sync|imem_rst), .re(imem_re), .wstrb(4'b0000),
           .a(imem_addr), .wd(32'd0),
           .rd(imem_data));

    mem #(DMEM_TYPE, SYNTH_DMEM_SIZE, BSRAM_DMEM_SIZE, DMEM_INIT_FILE) dmem
          (.clk(clk_dmem), .reset(rst_sync), .re(1'b1), .wstrb(dmem_Write),
           .a(dmem_Addr), .wd(dmem_WriteData),
           .rd(dmem_ReadData));
endmodule